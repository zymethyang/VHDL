`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:22:49 09/06/2018 
// Design Name: 
// Module Name:    GIAIMA_SELECT_INS_E 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module GIAIMA_SELECT_INS_E(
    input [2:0] I,
    output [7:0] O
    );


endmodule
